/* Copyright (C) 
* 
* This program is free software; you can redistribute it and/or
* modify it under the terms of the GNU General Public License
* as published by the Free Software Foundation; either version 2
* of the License, or (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program; if not, write to the Free Software
* Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  02111-1307, USA.
* 
* 2020 - Junying Hu
*/

package SimBench;

// ================================================================
// Modules Importation

// ================================================================
// Macro definition

// ================================================================
// Interface definition
//interface Multiplexer_IFC;
interface SimBench_IFC;
   method Action start;
   method ActionValue #(int) finish;
endinterface

// ================================================================
// Type Definition
typedef enum {IDLE, PROCESS, FINISH} State_MTB
deriving (Eq, Bits, FShow);

// ================================================================
// Module definition

endpackage
